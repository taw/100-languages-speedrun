module oddeven(A, O);
  input [15:0] A;
  output O;

  assign O = A[0];
endmodule
